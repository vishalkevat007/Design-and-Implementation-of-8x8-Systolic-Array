/scratch/asicfab/a/vkevat/systolic_design/LEF/gsclib045_tech.lef