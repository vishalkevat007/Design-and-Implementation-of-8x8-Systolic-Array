/scratch/asicfab/a/vkevat/systolic_design/LEF/gsclib045_macro.lef