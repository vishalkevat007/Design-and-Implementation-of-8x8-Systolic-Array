/scratch/asicfab/a/vkevat/Design-and-Implementation-of-8x8-Systolic-Array/LEF/gsclib045_tech.lef